module full_adder_4_bit (
    input  wire [3:0] a,
    input  wire [3:0] b,
    input  wire cin,
    output wire [3:0] sum,
    output wire cout
);
    // TODO: Implement the 4-bit full adder here
    assign {cout,sum} = a+b+cin;

endmodule
